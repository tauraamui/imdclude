module imdclude

pub fn backup_document(doc Document) ? {
	return error("backing up documents is not implemented")
}
